module NOT(b,a);
  input wire a;
  output wire b;
  
  assign b=~a;
endmodule
