module AND_2ip(c,a,b);
  input wire a,b;
  output wire c;
  
  assign c=a&b;
endmodule
